// Implement one cycle access by a voltage control: clk=0, precharge; clk=1, WL turn on
module bank_ctrl (

);

endmodule