module clk_copy (
    input clk,
    input clk_inv,
    input rst_n,
    output clk_copy
);

endmodule
